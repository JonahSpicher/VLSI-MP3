magic
tech sky130A
timestamp 1616551804
<< nwell >>
rect -180 705 2290 1710
rect 905 685 2290 705
<< nmos >>
rect -130 275 -80 575
rect -30 275 20 575
rect 70 275 120 575
rect 170 275 220 575
rect 270 275 320 575
rect 370 275 420 575
rect 470 275 520 575
rect 570 275 620 575
rect 670 275 720 575
rect 770 275 820 575
rect 970 275 1020 575
rect 1070 275 1120 575
rect 1250 275 1300 575
rect 1350 275 1400 575
rect 1530 275 1580 575
rect 1630 275 1680 575
rect 1810 275 1860 575
rect 1910 275 1960 575
rect 2090 275 2140 575
rect 2190 275 2240 575
<< pmos >>
rect 260 1315 310 1615
rect 360 1315 410 1615
rect 460 1315 510 1615
rect 560 1315 610 1615
rect 660 1315 710 1615
rect 760 1315 810 1615
rect 860 1315 910 1615
rect 960 1315 1010 1615
rect 1140 1315 1190 1615
rect 1240 1315 1290 1615
rect 1420 1315 1470 1615
rect 1520 1315 1570 1615
rect 1700 1315 1750 1615
rect 1800 1315 1850 1615
rect 1980 1315 2030 1615
rect 2080 1315 2130 1615
rect -45 785 5 1085
rect 55 785 105 1085
rect 155 785 205 1085
rect 255 785 305 1085
rect 355 785 405 1085
rect 455 785 505 1085
rect 555 785 605 1085
rect 655 785 705 1085
rect 755 785 805 1085
rect 855 785 905 1085
rect 1055 785 1105 1085
rect 1155 785 1205 1085
rect 1255 785 1305 1085
rect 1355 785 1405 1085
rect 1455 785 1505 1085
rect 1555 785 1605 1085
rect 1655 785 1705 1085
rect 1755 785 1805 1085
rect 1855 785 1905 1085
rect 1955 785 2005 1085
<< ndiff >>
rect -180 560 -130 575
rect -180 290 -165 560
rect -145 290 -130 560
rect -180 275 -130 290
rect -80 560 -30 575
rect -80 290 -65 560
rect -45 290 -30 560
rect -80 275 -30 290
rect 20 560 70 575
rect 20 290 35 560
rect 55 290 70 560
rect 20 275 70 290
rect 120 560 170 575
rect 120 290 135 560
rect 155 290 170 560
rect 120 275 170 290
rect 220 560 270 575
rect 220 290 235 560
rect 255 290 270 560
rect 220 275 270 290
rect 320 560 370 575
rect 320 290 335 560
rect 355 290 370 560
rect 320 275 370 290
rect 420 560 470 575
rect 420 290 435 560
rect 455 290 470 560
rect 420 275 470 290
rect 520 560 570 575
rect 520 290 535 560
rect 555 290 570 560
rect 520 275 570 290
rect 620 560 670 575
rect 620 290 635 560
rect 655 290 670 560
rect 620 275 670 290
rect 720 560 770 575
rect 720 290 735 560
rect 755 290 770 560
rect 720 275 770 290
rect 820 560 870 575
rect 920 560 970 575
rect 820 290 835 560
rect 855 290 870 560
rect 920 290 935 560
rect 955 290 970 560
rect 820 275 870 290
rect 920 275 970 290
rect 1020 560 1070 575
rect 1020 290 1035 560
rect 1055 290 1070 560
rect 1020 275 1070 290
rect 1120 560 1170 575
rect 1120 290 1135 560
rect 1155 290 1170 560
rect 1120 275 1170 290
rect 1200 560 1250 575
rect 1200 290 1215 560
rect 1235 290 1250 560
rect 1200 275 1250 290
rect 1300 560 1350 575
rect 1300 290 1315 560
rect 1335 290 1350 560
rect 1300 275 1350 290
rect 1400 560 1450 575
rect 1400 290 1415 560
rect 1435 290 1450 560
rect 1400 275 1450 290
rect 1480 560 1530 575
rect 1480 290 1495 560
rect 1515 290 1530 560
rect 1480 275 1530 290
rect 1580 560 1630 575
rect 1580 290 1595 560
rect 1615 290 1630 560
rect 1580 275 1630 290
rect 1680 560 1730 575
rect 1680 290 1695 560
rect 1715 290 1730 560
rect 1680 275 1730 290
rect 1760 560 1810 575
rect 1760 290 1775 560
rect 1795 290 1810 560
rect 1760 275 1810 290
rect 1860 560 1910 575
rect 1860 290 1875 560
rect 1895 290 1910 560
rect 1860 275 1910 290
rect 1960 560 2010 575
rect 1960 290 1975 560
rect 1995 290 2010 560
rect 1960 275 2010 290
rect 2040 560 2090 575
rect 2040 290 2055 560
rect 2075 290 2090 560
rect 2040 275 2090 290
rect 2140 560 2190 575
rect 2140 290 2155 560
rect 2175 290 2190 560
rect 2140 275 2190 290
rect 2240 560 2290 575
rect 2240 290 2255 560
rect 2275 290 2290 560
rect 2240 275 2290 290
<< pdiff >>
rect 210 1600 260 1615
rect 210 1330 225 1600
rect 245 1330 260 1600
rect 210 1315 260 1330
rect 310 1600 360 1615
rect 310 1330 325 1600
rect 345 1330 360 1600
rect 310 1315 360 1330
rect 410 1600 460 1615
rect 410 1330 425 1600
rect 445 1330 460 1600
rect 410 1315 460 1330
rect 510 1600 560 1615
rect 510 1330 525 1600
rect 545 1330 560 1600
rect 510 1315 560 1330
rect 610 1600 660 1615
rect 610 1330 625 1600
rect 645 1330 660 1600
rect 610 1315 660 1330
rect 710 1600 760 1615
rect 710 1330 725 1600
rect 745 1330 760 1600
rect 710 1315 760 1330
rect 810 1600 860 1615
rect 810 1330 825 1600
rect 845 1330 860 1600
rect 810 1315 860 1330
rect 910 1600 960 1615
rect 910 1330 925 1600
rect 945 1330 960 1600
rect 910 1315 960 1330
rect 1010 1600 1060 1615
rect 1010 1330 1025 1600
rect 1045 1330 1060 1600
rect 1010 1315 1060 1330
rect 1090 1600 1140 1615
rect 1090 1330 1105 1600
rect 1125 1330 1140 1600
rect 1090 1315 1140 1330
rect 1190 1600 1240 1615
rect 1190 1330 1205 1600
rect 1225 1330 1240 1600
rect 1190 1315 1240 1330
rect 1290 1600 1340 1615
rect 1290 1330 1305 1600
rect 1325 1330 1340 1600
rect 1290 1315 1340 1330
rect 1370 1600 1420 1615
rect 1370 1330 1385 1600
rect 1405 1330 1420 1600
rect 1370 1315 1420 1330
rect 1470 1600 1520 1615
rect 1470 1330 1485 1600
rect 1505 1330 1520 1600
rect 1470 1315 1520 1330
rect 1570 1600 1620 1615
rect 1570 1330 1585 1600
rect 1605 1330 1620 1600
rect 1570 1315 1620 1330
rect 1650 1600 1700 1615
rect 1650 1330 1665 1600
rect 1685 1330 1700 1600
rect 1650 1315 1700 1330
rect 1750 1600 1800 1615
rect 1750 1330 1765 1600
rect 1785 1330 1800 1600
rect 1750 1315 1800 1330
rect 1850 1600 1900 1615
rect 1850 1330 1865 1600
rect 1885 1330 1900 1600
rect 1850 1315 1900 1330
rect 1930 1600 1980 1615
rect 1930 1330 1945 1600
rect 1965 1330 1980 1600
rect 1930 1315 1980 1330
rect 2030 1600 2080 1615
rect 2030 1330 2045 1600
rect 2065 1330 2080 1600
rect 2030 1315 2080 1330
rect 2130 1600 2180 1615
rect 2130 1330 2145 1600
rect 2165 1330 2180 1600
rect 2130 1315 2180 1330
rect -95 1070 -45 1085
rect -95 800 -80 1070
rect -60 800 -45 1070
rect -95 785 -45 800
rect 5 1070 55 1085
rect 5 800 20 1070
rect 40 800 55 1070
rect 5 785 55 800
rect 105 1070 155 1085
rect 105 800 120 1070
rect 140 800 155 1070
rect 105 785 155 800
rect 205 1070 255 1085
rect 205 800 220 1070
rect 240 800 255 1070
rect 205 785 255 800
rect 305 1070 355 1085
rect 305 800 320 1070
rect 340 800 355 1070
rect 305 785 355 800
rect 405 1070 455 1085
rect 405 800 420 1070
rect 440 800 455 1070
rect 405 785 455 800
rect 505 1070 555 1085
rect 505 800 520 1070
rect 540 800 555 1070
rect 505 785 555 800
rect 605 1070 655 1085
rect 605 800 620 1070
rect 640 800 655 1070
rect 605 785 655 800
rect 705 1070 755 1085
rect 705 800 720 1070
rect 740 800 755 1070
rect 705 785 755 800
rect 805 1070 855 1085
rect 805 800 820 1070
rect 840 800 855 1070
rect 805 785 855 800
rect 905 1070 955 1085
rect 1005 1070 1055 1085
rect 905 800 920 1070
rect 940 800 955 1070
rect 1005 800 1020 1070
rect 1040 800 1055 1070
rect 905 785 955 800
rect 1005 785 1055 800
rect 1105 1070 1155 1085
rect 1105 800 1120 1070
rect 1140 800 1155 1070
rect 1105 785 1155 800
rect 1205 1070 1255 1085
rect 1205 800 1220 1070
rect 1240 800 1255 1070
rect 1205 785 1255 800
rect 1305 1070 1355 1085
rect 1305 800 1320 1070
rect 1340 800 1355 1070
rect 1305 785 1355 800
rect 1405 1070 1455 1085
rect 1405 800 1420 1070
rect 1440 800 1455 1070
rect 1405 785 1455 800
rect 1505 1070 1555 1085
rect 1505 800 1520 1070
rect 1540 800 1555 1070
rect 1505 785 1555 800
rect 1605 1070 1655 1085
rect 1605 800 1620 1070
rect 1640 800 1655 1070
rect 1605 785 1655 800
rect 1705 1070 1755 1085
rect 1705 800 1720 1070
rect 1740 800 1755 1070
rect 1705 785 1755 800
rect 1805 1070 1855 1085
rect 1805 800 1820 1070
rect 1840 800 1855 1070
rect 1805 785 1855 800
rect 1905 1070 1955 1085
rect 1905 800 1920 1070
rect 1940 800 1955 1070
rect 1905 785 1955 800
rect 2005 1070 2055 1085
rect 2005 800 2020 1070
rect 2040 800 2055 1070
rect 2005 785 2055 800
<< ndiffc >>
rect -165 290 -145 560
rect -65 290 -45 560
rect 35 290 55 560
rect 135 290 155 560
rect 235 290 255 560
rect 335 290 355 560
rect 435 290 455 560
rect 535 290 555 560
rect 635 290 655 560
rect 735 290 755 560
rect 835 290 855 560
rect 935 290 955 560
rect 1035 290 1055 560
rect 1135 290 1155 560
rect 1215 290 1235 560
rect 1315 290 1335 560
rect 1415 290 1435 560
rect 1495 290 1515 560
rect 1595 290 1615 560
rect 1695 290 1715 560
rect 1775 290 1795 560
rect 1875 290 1895 560
rect 1975 290 1995 560
rect 2055 290 2075 560
rect 2155 290 2175 560
rect 2255 290 2275 560
<< pdiffc >>
rect 225 1330 245 1600
rect 325 1330 345 1600
rect 425 1330 445 1600
rect 525 1330 545 1600
rect 625 1330 645 1600
rect 725 1330 745 1600
rect 825 1330 845 1600
rect 925 1330 945 1600
rect 1025 1330 1045 1600
rect 1105 1330 1125 1600
rect 1205 1330 1225 1600
rect 1305 1330 1325 1600
rect 1385 1330 1405 1600
rect 1485 1330 1505 1600
rect 1585 1330 1605 1600
rect 1665 1330 1685 1600
rect 1765 1330 1785 1600
rect 1865 1330 1885 1600
rect 1945 1330 1965 1600
rect 2045 1330 2065 1600
rect 2145 1330 2165 1600
rect -80 800 -60 1070
rect 20 800 40 1070
rect 120 800 140 1070
rect 220 800 240 1070
rect 320 800 340 1070
rect 420 800 440 1070
rect 520 800 540 1070
rect 620 800 640 1070
rect 720 800 740 1070
rect 820 800 840 1070
rect 920 800 940 1070
rect 1020 800 1040 1070
rect 1120 800 1140 1070
rect 1220 800 1240 1070
rect 1320 800 1340 1070
rect 1420 800 1440 1070
rect 1520 800 1540 1070
rect 1620 800 1640 1070
rect 1720 800 1740 1070
rect 1820 800 1840 1070
rect 1920 800 1940 1070
rect 2020 800 2040 1070
<< psubdiff >>
rect 870 560 920 575
rect 870 290 885 560
rect 905 290 920 560
rect 870 275 920 290
<< nsubdiff >>
rect 160 1600 210 1615
rect 160 1330 175 1600
rect 195 1330 210 1600
rect 160 1315 210 1330
rect 955 1070 1005 1085
rect 955 800 970 1070
rect 990 800 1005 1070
rect 955 785 1005 800
<< psubdiffcont >>
rect 885 290 905 560
<< nsubdiffcont >>
rect 175 1330 195 1600
rect 970 800 990 1070
<< poly >>
rect 2015 1700 2055 1710
rect 2015 1680 2025 1700
rect 2045 1680 2055 1700
rect 260 1660 300 1670
rect 260 1640 270 1660
rect 290 1640 300 1660
rect 2015 1655 2055 1680
rect 2015 1640 2030 1655
rect 260 1630 300 1640
rect 260 1615 310 1630
rect 360 1625 710 1640
rect 360 1615 410 1625
rect 460 1615 510 1625
rect 560 1615 610 1625
rect 660 1615 710 1625
rect 760 1615 810 1630
rect 860 1615 910 1630
rect 960 1625 2030 1640
rect 960 1615 1010 1625
rect 1140 1615 1190 1625
rect 1240 1615 1290 1625
rect 1420 1615 1470 1625
rect 1520 1615 1570 1625
rect 1700 1615 1750 1625
rect 1800 1615 1850 1625
rect 1980 1615 2030 1625
rect 2080 1615 2130 1630
rect 260 1300 310 1315
rect 360 1300 410 1315
rect 460 1300 510 1315
rect 560 1300 610 1315
rect 660 1300 710 1315
rect 760 1305 810 1315
rect 860 1305 910 1315
rect 760 1300 910 1305
rect 960 1300 1010 1315
rect 1140 1300 1190 1315
rect 1240 1300 1290 1315
rect 1420 1300 1470 1315
rect 1520 1300 1570 1315
rect 1700 1300 1750 1315
rect 1800 1300 1850 1315
rect 1980 1300 2030 1315
rect 2080 1300 2130 1315
rect 360 1290 400 1300
rect 795 1290 880 1300
rect 360 1270 370 1290
rect 390 1270 400 1290
rect 360 1260 400 1270
rect 65 1155 105 1165
rect -45 1130 -5 1140
rect -45 1110 -35 1130
rect -15 1110 -5 1130
rect 65 1135 75 1155
rect 95 1140 105 1155
rect 865 1140 880 1290
rect 2090 1290 2130 1300
rect 2090 1270 2100 1290
rect 2120 1270 2130 1290
rect 2090 1260 2130 1270
rect 1855 1250 1895 1260
rect 1855 1230 1865 1250
rect 1885 1230 1895 1250
rect 1855 1220 1895 1230
rect 95 1135 770 1140
rect 65 1125 770 1135
rect -45 1100 -5 1110
rect 90 1100 105 1125
rect 390 1100 405 1125
rect -45 1085 5 1100
rect 55 1085 105 1100
rect 155 1085 205 1100
rect 255 1085 305 1100
rect 355 1085 405 1100
rect 455 1100 470 1125
rect 755 1100 770 1125
rect 865 1130 905 1140
rect 865 1110 875 1130
rect 895 1110 905 1130
rect 865 1100 905 1110
rect 455 1085 505 1100
rect 555 1085 605 1100
rect 655 1085 705 1100
rect 755 1085 805 1100
rect 855 1085 905 1100
rect 1055 1130 1095 1140
rect 1055 1110 1065 1130
rect 1085 1110 1095 1130
rect 1055 1100 1095 1110
rect 1855 1100 1875 1220
rect 1965 1130 2005 1140
rect 1965 1110 1975 1130
rect 1995 1110 2005 1130
rect 1965 1100 2005 1110
rect 1055 1085 1105 1100
rect 1155 1085 1205 1100
rect 1255 1085 1305 1100
rect 1355 1085 1405 1100
rect 1455 1085 1505 1100
rect 1555 1085 1605 1100
rect 1655 1085 1705 1100
rect 1755 1085 1805 1100
rect 1855 1085 1905 1100
rect 1955 1085 2005 1100
rect -45 770 5 785
rect 55 770 105 785
rect 155 770 205 785
rect 255 770 305 785
rect 355 770 405 785
rect 455 770 505 785
rect 555 770 605 785
rect 655 770 705 785
rect 755 770 805 785
rect 855 770 905 785
rect 1055 770 1105 785
rect 1155 775 1205 785
rect 1255 775 1305 785
rect 1355 775 1405 785
rect 1455 775 1505 785
rect 1555 775 1605 785
rect 1655 775 1705 785
rect 1755 775 1805 785
rect 1855 775 1905 785
rect 155 755 270 770
rect 155 745 170 755
rect -180 735 170 745
rect -180 715 -170 735
rect -150 730 170 735
rect 255 745 270 755
rect 590 755 670 770
rect 1155 760 1905 775
rect 1955 770 2005 785
rect 590 745 605 755
rect 255 730 605 745
rect 1705 740 1715 760
rect 1735 740 1745 760
rect 1705 730 1745 740
rect -150 715 -140 730
rect -180 705 -140 715
rect 2250 680 2290 690
rect -180 670 -140 680
rect -180 650 -170 670
rect -150 655 -15 670
rect -150 650 -140 655
rect -180 640 -140 650
rect -120 620 -80 630
rect -120 600 -110 620
rect -90 600 -80 620
rect -120 590 -80 600
rect -130 575 -80 590
rect -30 600 -15 655
rect 210 660 250 670
rect 210 640 220 660
rect 240 645 250 660
rect 575 660 615 670
rect 2250 665 2260 680
rect 575 645 585 660
rect 240 640 585 645
rect 605 640 615 660
rect 210 630 615 640
rect 1145 655 1285 665
rect 1145 635 1155 655
rect 1175 650 1255 655
rect 1175 635 1185 650
rect 1145 625 1185 635
rect 1245 635 1255 650
rect 1275 635 1285 655
rect 1245 625 1285 635
rect 2125 660 2260 665
rect 2280 660 2290 680
rect 2125 650 2290 660
rect 780 615 820 625
rect -30 585 720 600
rect 780 595 790 615
rect 810 595 820 615
rect 780 590 820 595
rect -30 575 20 585
rect 70 575 120 585
rect 170 575 220 585
rect 270 575 320 585
rect 370 575 420 585
rect 470 575 520 585
rect 570 575 620 585
rect 670 575 720 585
rect 770 575 820 590
rect 970 615 1010 625
rect 970 595 980 615
rect 1000 595 1010 615
rect 2125 600 2140 650
rect 970 590 1010 595
rect 970 575 1020 590
rect 1070 585 2140 600
rect 2200 615 2240 625
rect 2200 595 2210 615
rect 2230 595 2240 615
rect 2200 590 2240 595
rect 1070 575 1120 585
rect 1250 575 1300 585
rect 1350 575 1400 585
rect 1530 575 1580 585
rect 1630 575 1680 585
rect 1810 575 1860 585
rect 1910 575 1960 585
rect 2090 575 2140 585
rect 2190 575 2240 590
rect -130 260 -80 275
rect -30 260 20 275
rect 70 260 120 275
rect 170 260 220 275
rect 270 260 320 275
rect 370 260 420 275
rect 470 260 520 275
rect 570 260 620 275
rect 670 260 720 275
rect 770 260 820 275
rect 970 260 1020 275
rect 1070 260 1120 275
rect 1250 260 1300 275
rect 1350 260 1400 275
rect 1425 255 1465 265
rect 1530 260 1580 275
rect 1630 260 1680 275
rect 1425 235 1435 255
rect 1455 235 1465 255
rect 1745 255 1785 265
rect 1810 260 1860 275
rect 1910 260 1960 275
rect 2090 260 2140 275
rect 2190 260 2240 275
rect 1745 235 1755 255
rect 1775 235 1785 255
rect 1425 220 1785 235
<< polycont >>
rect 2025 1680 2045 1700
rect 270 1640 290 1660
rect 370 1270 390 1290
rect -35 1110 -15 1130
rect 75 1135 95 1155
rect 2100 1270 2120 1290
rect 1865 1230 1885 1250
rect 875 1110 895 1130
rect 1065 1110 1085 1130
rect 1975 1110 1995 1130
rect -170 715 -150 735
rect 1715 740 1735 760
rect -170 650 -150 670
rect -110 600 -90 620
rect 220 640 240 660
rect 585 640 605 660
rect 1155 635 1175 655
rect 1255 635 1275 655
rect 2260 660 2280 680
rect 790 595 810 615
rect 980 595 1000 615
rect 2210 595 2230 615
rect 1435 235 1455 255
rect 1755 235 1775 255
<< locali >>
rect 1115 1690 1875 1710
rect 260 1660 300 1670
rect 260 1650 270 1660
rect 235 1640 270 1650
rect 290 1640 300 1660
rect 235 1630 300 1640
rect 335 1630 735 1650
rect 235 1610 255 1630
rect 335 1610 355 1630
rect 525 1610 545 1630
rect 715 1610 735 1630
rect 1115 1610 1135 1690
rect 1215 1660 1290 1670
rect 1215 1640 1225 1660
rect 1280 1640 1290 1660
rect 1215 1630 1290 1640
rect 1215 1610 1235 1630
rect 1315 1610 1335 1690
rect 1655 1610 1675 1690
rect 1700 1660 1775 1670
rect 1700 1640 1710 1660
rect 1765 1640 1775 1660
rect 1700 1630 1775 1640
rect 1755 1610 1775 1630
rect 1855 1650 1875 1690
rect 2015 1700 2055 1710
rect 2015 1680 2025 1700
rect 2045 1680 2055 1700
rect 2015 1670 2055 1680
rect 1855 1630 2235 1650
rect 1855 1610 1875 1630
rect 165 1600 255 1610
rect 165 1330 175 1600
rect 195 1330 225 1600
rect 245 1330 255 1600
rect 165 1320 255 1330
rect 315 1600 355 1610
rect 315 1330 325 1600
rect 345 1330 355 1600
rect 315 1320 355 1330
rect 415 1600 455 1610
rect 415 1330 425 1600
rect 445 1330 455 1600
rect 415 1320 455 1330
rect 515 1600 555 1610
rect 515 1330 525 1600
rect 545 1330 555 1600
rect 515 1320 555 1330
rect 615 1600 655 1610
rect 615 1330 625 1600
rect 645 1330 655 1600
rect 615 1320 655 1330
rect 715 1600 755 1610
rect 715 1330 725 1600
rect 745 1330 755 1600
rect 715 1320 755 1330
rect 815 1600 855 1610
rect 815 1330 825 1600
rect 845 1330 855 1600
rect 815 1320 855 1330
rect 915 1600 955 1610
rect 915 1330 925 1600
rect 945 1330 955 1600
rect 915 1320 955 1330
rect 1015 1600 1055 1610
rect 1015 1330 1025 1600
rect 1045 1330 1055 1600
rect 1015 1320 1055 1330
rect 1095 1600 1135 1610
rect 1095 1330 1105 1600
rect 1125 1330 1135 1600
rect 1095 1320 1135 1330
rect 1195 1600 1235 1610
rect 1195 1330 1205 1600
rect 1225 1330 1235 1600
rect 1195 1320 1235 1330
rect 1295 1600 1335 1610
rect 1295 1330 1305 1600
rect 1325 1330 1335 1600
rect 1295 1320 1335 1330
rect 1375 1600 1415 1610
rect 1375 1330 1385 1600
rect 1405 1330 1415 1600
rect 1375 1320 1415 1330
rect 1475 1600 1515 1610
rect 1475 1330 1485 1600
rect 1505 1330 1515 1600
rect 1475 1320 1515 1330
rect 1575 1600 1615 1610
rect 1575 1330 1585 1600
rect 1605 1330 1615 1600
rect 1575 1320 1615 1330
rect 1655 1600 1695 1610
rect 1655 1330 1665 1600
rect 1685 1330 1695 1600
rect 1655 1320 1695 1330
rect 1755 1600 1795 1610
rect 1755 1330 1765 1600
rect 1785 1330 1795 1600
rect 1755 1320 1795 1330
rect 1855 1600 1895 1610
rect 1855 1330 1865 1600
rect 1885 1330 1895 1600
rect 1855 1320 1895 1330
rect 1935 1600 1975 1610
rect 1935 1330 1945 1600
rect 1965 1330 1975 1600
rect 1935 1320 1975 1330
rect 2035 1600 2075 1610
rect 2035 1330 2045 1600
rect 2065 1330 2075 1600
rect 2035 1320 2075 1330
rect 2135 1600 2175 1610
rect 2135 1330 2145 1600
rect 2165 1330 2175 1600
rect 2135 1320 2175 1330
rect -180 1295 145 1315
rect 125 1280 145 1295
rect 360 1290 400 1300
rect 360 1280 370 1290
rect 125 1270 370 1280
rect 390 1270 400 1290
rect 125 1260 400 1270
rect 535 1280 555 1320
rect 535 1260 650 1280
rect -180 1190 -105 1200
rect -180 1170 -170 1190
rect -115 1180 -105 1190
rect -115 1170 105 1180
rect -180 1160 105 1170
rect 65 1155 105 1160
rect -45 1130 -5 1140
rect -45 1120 -35 1130
rect -70 1110 -35 1120
rect -15 1110 -5 1130
rect 65 1135 75 1155
rect 95 1135 105 1155
rect 65 1125 105 1135
rect 630 1120 650 1260
rect 935 1240 955 1320
rect 1035 1300 1055 1320
rect 1375 1300 1395 1320
rect 1035 1290 1450 1300
rect 1035 1280 1385 1290
rect 1375 1270 1385 1280
rect 1440 1270 1450 1290
rect 1375 1260 1450 1270
rect 1485 1240 1505 1320
rect 1595 1300 1615 1320
rect 1935 1300 1955 1320
rect 1540 1290 1955 1300
rect 1540 1270 1550 1290
rect 1605 1280 1955 1290
rect 1605 1270 1615 1280
rect 1540 1260 1615 1270
rect 1855 1250 1895 1260
rect 1855 1240 1865 1250
rect 935 1230 1865 1240
rect 1885 1240 1895 1250
rect 2035 1240 2055 1320
rect 2135 1300 2155 1320
rect 2090 1290 2155 1300
rect 2090 1270 2100 1290
rect 2120 1280 2155 1290
rect 2120 1270 2130 1280
rect 2090 1260 2130 1270
rect 1885 1230 2055 1240
rect 935 1220 2055 1230
rect 1575 1190 1650 1200
rect 1575 1180 1585 1190
rect 1130 1170 1585 1180
rect 1640 1180 1650 1190
rect 1640 1170 1930 1180
rect 1130 1160 1930 1170
rect 865 1130 905 1140
rect -70 1100 -5 1110
rect 130 1100 730 1120
rect 865 1110 875 1130
rect 895 1120 905 1130
rect 1055 1130 1095 1140
rect 1055 1120 1065 1130
rect 895 1110 950 1120
rect 865 1100 950 1110
rect -70 1080 -50 1100
rect 130 1080 150 1100
rect 330 1080 350 1100
rect 510 1080 530 1100
rect 710 1080 730 1100
rect 930 1080 950 1100
rect 1030 1110 1065 1120
rect 1085 1110 1095 1130
rect 1030 1100 1095 1110
rect 1030 1080 1050 1100
rect 1130 1080 1150 1160
rect 1310 1130 1385 1140
rect 1310 1110 1320 1130
rect 1375 1110 1385 1130
rect 1310 1100 1385 1110
rect 1310 1080 1330 1100
rect 1520 1080 1540 1160
rect 1675 1130 1750 1140
rect 1675 1110 1685 1130
rect 1740 1110 1750 1130
rect 1675 1100 1750 1110
rect 1730 1080 1750 1100
rect 1910 1080 1930 1160
rect 1965 1130 2005 1140
rect 1965 1110 1975 1130
rect 1995 1120 2005 1130
rect 1995 1110 2030 1120
rect 1965 1100 2030 1110
rect 2010 1080 2030 1100
rect -90 1070 -50 1080
rect -90 800 -80 1070
rect -60 800 -50 1070
rect -90 790 -50 800
rect 10 1070 50 1080
rect 10 800 20 1070
rect 40 800 50 1070
rect 10 790 50 800
rect 110 1070 150 1080
rect 110 800 120 1070
rect 140 800 150 1070
rect 110 790 150 800
rect 210 1070 250 1080
rect 210 800 220 1070
rect 240 800 250 1070
rect 210 790 250 800
rect 310 1070 350 1080
rect 310 800 320 1070
rect 340 800 350 1070
rect 310 790 350 800
rect 410 1070 450 1080
rect 410 800 420 1070
rect 440 800 450 1070
rect 410 790 450 800
rect 510 1070 550 1080
rect 510 800 520 1070
rect 540 800 550 1070
rect 510 790 550 800
rect 610 1070 650 1080
rect 610 800 620 1070
rect 640 800 650 1070
rect 610 790 650 800
rect 710 1070 750 1080
rect 710 800 720 1070
rect 740 800 750 1070
rect 710 790 750 800
rect 810 1070 850 1080
rect 810 800 820 1070
rect 840 800 850 1070
rect 810 790 850 800
rect 910 1070 1050 1080
rect 910 800 920 1070
rect 940 800 970 1070
rect 990 800 1020 1070
rect 1040 800 1050 1070
rect 910 790 1050 800
rect 1110 1070 1150 1080
rect 1110 800 1120 1070
rect 1140 800 1150 1070
rect 1110 790 1150 800
rect 1210 1070 1250 1080
rect 1210 800 1220 1070
rect 1240 800 1250 1070
rect 1210 790 1250 800
rect 1310 1070 1350 1080
rect 1310 800 1320 1070
rect 1340 800 1350 1070
rect 1310 790 1350 800
rect 1410 1070 1450 1080
rect 1410 800 1420 1070
rect 1440 800 1450 1070
rect 1410 790 1450 800
rect 1510 1070 1550 1080
rect 1510 800 1520 1070
rect 1540 800 1550 1070
rect 1510 790 1550 800
rect 1610 1070 1650 1080
rect 1610 800 1620 1070
rect 1640 800 1650 1070
rect 1610 790 1650 800
rect 1710 1070 1750 1080
rect 1710 800 1720 1070
rect 1740 800 1750 1070
rect 1710 790 1750 800
rect 1810 1070 1850 1080
rect 1810 800 1820 1070
rect 1840 800 1850 1070
rect 1810 790 1850 800
rect 1910 1070 1950 1080
rect 1910 800 1920 1070
rect 1940 800 1950 1070
rect 1910 790 1950 800
rect 2010 1070 2050 1080
rect 2010 800 2020 1070
rect 2040 800 2050 1070
rect 2010 790 2050 800
rect -180 735 -105 745
rect -180 715 -170 735
rect -115 715 -105 735
rect -180 705 -105 715
rect 30 710 50 790
rect 210 770 230 790
rect 210 760 285 770
rect 210 740 220 760
rect 275 740 285 760
rect 210 730 285 740
rect 430 710 450 790
rect 630 770 650 790
rect 575 760 650 770
rect 575 740 585 760
rect 640 740 650 760
rect 575 730 650 740
rect 810 710 830 790
rect 30 690 830 710
rect 1705 760 1745 770
rect 2215 765 2235 1630
rect 1705 740 1715 760
rect 1735 740 1745 760
rect 1705 730 1745 740
rect 2160 755 2235 765
rect 2160 735 2170 755
rect 2225 735 2235 755
rect -180 670 -140 680
rect -180 650 -170 670
rect -150 650 -140 670
rect 210 660 250 670
rect 210 650 220 660
rect -180 640 -140 650
rect 145 640 220 650
rect 240 640 250 660
rect 145 630 250 640
rect -120 620 -80 630
rect -120 610 -110 620
rect -155 600 -110 610
rect -90 600 -80 620
rect -155 590 -80 600
rect -155 570 -135 590
rect 145 570 165 630
rect 345 570 365 690
rect 905 685 1225 705
rect 905 670 925 685
rect 575 660 925 670
rect 575 650 585 660
rect 545 640 585 650
rect 640 650 925 660
rect 1145 655 1185 665
rect 640 640 650 650
rect 545 630 650 640
rect 1145 635 1155 655
rect 1175 635 1185 655
rect 545 570 565 630
rect 1145 625 1185 635
rect 780 615 820 625
rect 780 595 790 615
rect 810 605 820 615
rect 970 615 1010 625
rect 970 605 980 615
rect 810 595 845 605
rect 780 585 845 595
rect 825 570 845 585
rect 945 595 980 605
rect 1000 595 1010 615
rect 945 585 1010 595
rect 945 570 965 585
rect 1145 570 1165 625
rect -180 560 -135 570
rect -180 290 -165 560
rect -145 290 -135 560
rect -180 280 -135 290
rect -75 560 -35 570
rect -75 290 -65 560
rect -45 290 -35 560
rect -75 280 -35 290
rect 25 560 65 570
rect 25 290 35 560
rect 55 290 65 560
rect 25 280 65 290
rect 125 560 165 570
rect 125 290 135 560
rect 155 290 165 560
rect 125 280 165 290
rect 225 560 265 570
rect 225 290 235 560
rect 255 290 265 560
rect 225 280 265 290
rect 325 560 365 570
rect 325 290 335 560
rect 355 290 365 560
rect 325 280 365 290
rect 425 560 465 570
rect 425 290 435 560
rect 455 290 465 560
rect 425 280 465 290
rect 525 560 565 570
rect 525 290 535 560
rect 555 290 565 560
rect 525 280 565 290
rect 625 560 665 570
rect 625 290 635 560
rect 655 290 665 560
rect 625 280 665 290
rect 725 560 765 570
rect 725 290 735 560
rect 755 290 765 560
rect 725 280 765 290
rect 825 560 965 570
rect 825 290 835 560
rect 855 290 885 560
rect 905 290 935 560
rect 955 290 965 560
rect 825 280 965 290
rect 1025 560 1065 570
rect 1025 290 1035 560
rect 1055 290 1065 560
rect -55 255 -35 280
rect 345 255 365 280
rect 745 255 765 280
rect 1025 265 1065 290
rect 1125 560 1165 570
rect 1125 290 1135 560
rect 1155 290 1165 560
rect 1125 280 1165 290
rect 1205 570 1225 685
rect 1705 670 1725 730
rect 2160 725 2235 735
rect 2250 680 2290 690
rect 1245 655 2065 670
rect 1245 635 1255 655
rect 1275 650 2065 655
rect 2250 660 2260 680
rect 2280 660 2290 680
rect 2250 650 2290 660
rect 1275 635 1285 650
rect 1245 625 1285 635
rect 1325 620 1400 630
rect 1325 600 1335 620
rect 1390 600 1400 620
rect 1325 590 1400 600
rect 1325 570 1345 590
rect 1485 570 1505 650
rect 1705 570 1725 650
rect 1810 620 1885 630
rect 1810 600 1820 620
rect 1875 600 1885 620
rect 1810 590 1885 600
rect 1865 570 1885 590
rect 2045 570 2065 650
rect 2200 615 2240 625
rect 2200 595 2210 615
rect 2230 605 2240 615
rect 2230 595 2265 605
rect 2200 585 2265 595
rect 2245 570 2265 585
rect 1205 560 1245 570
rect 1205 290 1215 560
rect 1235 290 1245 560
rect 1205 280 1245 290
rect 1305 560 1345 570
rect 1305 290 1315 560
rect 1335 290 1345 560
rect 1305 280 1345 290
rect 1405 560 1445 570
rect 1405 290 1415 560
rect 1435 290 1445 560
rect 1405 280 1445 290
rect 1485 560 1525 570
rect 1485 290 1495 560
rect 1515 290 1525 560
rect 1485 280 1525 290
rect 1585 560 1625 570
rect 1585 290 1595 560
rect 1615 290 1625 560
rect 1025 255 1100 265
rect -55 235 1035 255
rect 1090 235 1100 255
rect 1025 225 1100 235
rect 1225 250 1245 280
rect 1425 265 1445 280
rect 1585 265 1625 290
rect 1685 560 1725 570
rect 1685 290 1695 560
rect 1715 290 1725 560
rect 1685 280 1725 290
rect 1765 560 1805 570
rect 1765 290 1775 560
rect 1795 290 1805 560
rect 1765 280 1805 290
rect 1865 560 1905 570
rect 1865 290 1875 560
rect 1895 290 1905 560
rect 1865 280 1905 290
rect 1965 560 2005 570
rect 1965 290 1975 560
rect 1995 290 2005 560
rect 1965 280 2005 290
rect 2045 560 2085 570
rect 2045 290 2055 560
rect 2075 290 2085 560
rect 2045 280 2085 290
rect 2145 560 2185 570
rect 2145 290 2155 560
rect 2175 290 2185 560
rect 1765 265 1785 280
rect 1425 255 1465 265
rect 1425 250 1435 255
rect 1225 235 1435 250
rect 1455 235 1465 255
rect 1225 230 1465 235
rect 1425 225 1465 230
rect 1585 255 1660 265
rect 1585 235 1595 255
rect 1650 235 1660 255
rect 1585 225 1660 235
rect 1745 255 1785 265
rect 1745 235 1755 255
rect 1775 250 1785 255
rect 1985 250 2005 280
rect 2145 265 2185 290
rect 2245 560 2285 570
rect 2245 290 2255 560
rect 2275 290 2285 560
rect 2245 280 2285 290
rect 1775 235 2005 250
rect 1745 230 2005 235
rect 2110 255 2185 265
rect 2110 235 2120 255
rect 2175 235 2185 255
rect 1745 225 1785 230
rect 2110 225 2185 235
<< viali >>
rect 1225 1640 1280 1660
rect 1710 1640 1765 1660
rect 175 1330 195 1600
rect 225 1330 245 1600
rect 425 1330 445 1600
rect 625 1330 645 1600
rect 825 1330 845 1600
rect 2145 1330 2165 1600
rect -170 1170 -115 1190
rect 1385 1270 1440 1290
rect 1550 1270 1605 1290
rect 1585 1170 1640 1190
rect 1320 1110 1375 1130
rect 1685 1110 1740 1130
rect -80 800 -60 1070
rect 920 800 940 1070
rect 970 800 990 1070
rect 1020 800 1040 1070
rect 1220 800 1240 1070
rect 1420 800 1440 1070
rect 1620 800 1640 1070
rect 1820 800 1840 1070
rect 2020 800 2040 1070
rect -170 715 -150 735
rect -150 715 -115 735
rect 220 740 275 760
rect 585 740 640 760
rect 2170 735 2225 755
rect 585 640 605 660
rect 605 640 640 660
rect -165 290 -145 560
rect 35 290 55 560
rect 235 290 255 560
rect 435 290 455 560
rect 635 290 655 560
rect 835 290 855 560
rect 885 290 905 560
rect 935 290 955 560
rect 1335 600 1390 620
rect 1820 600 1875 620
rect 1035 235 1090 255
rect 1595 235 1650 255
rect 2255 290 2275 560
rect 2120 235 2175 255
<< metal1 >>
rect 1215 1660 1775 1670
rect 1215 1640 1225 1660
rect 1280 1640 1710 1660
rect 1765 1640 1775 1660
rect 1215 1630 1775 1640
rect -180 1600 855 1610
rect -180 1330 175 1600
rect 195 1330 225 1600
rect 245 1330 425 1600
rect 445 1330 625 1600
rect 645 1330 825 1600
rect 845 1330 855 1600
rect -180 1320 855 1330
rect -180 1190 -105 1200
rect -180 1170 -170 1190
rect -115 1170 -105 1190
rect -180 1160 -105 1170
rect 815 1080 855 1320
rect 1375 1290 1615 1300
rect 1375 1270 1385 1290
rect 1440 1270 1550 1290
rect 1605 1270 1615 1290
rect 1375 1260 1615 1270
rect 1575 1200 1615 1260
rect 1575 1190 1650 1200
rect 1575 1170 1585 1190
rect 1640 1170 1650 1190
rect 1575 1160 1650 1170
rect 1675 1140 1695 1630
rect 2010 1600 2290 1610
rect 2010 1330 2145 1600
rect 2165 1330 2290 1600
rect 2010 1320 2290 1330
rect 1310 1130 1750 1140
rect 1310 1110 1320 1130
rect 1375 1110 1685 1130
rect 1740 1110 1750 1130
rect 1310 1100 1750 1110
rect 2010 1080 2050 1320
rect -90 1070 2290 1080
rect -90 800 -80 1070
rect -60 800 920 1070
rect 940 800 970 1070
rect 990 800 1020 1070
rect 1040 800 1220 1070
rect 1240 800 1420 1070
rect 1440 800 1620 1070
rect 1640 800 1820 1070
rect 1840 800 2020 1070
rect 2040 800 2290 1070
rect -90 790 2290 800
rect 210 760 650 770
rect -180 735 -105 745
rect -180 715 -170 735
rect -115 715 -105 735
rect 210 740 220 760
rect 275 740 585 760
rect 640 740 650 760
rect 210 730 650 740
rect -180 705 -105 715
rect 575 660 650 730
rect 575 640 585 660
rect 640 640 650 660
rect 575 630 650 640
rect 2115 755 2290 765
rect 2115 735 2170 755
rect 2225 735 2290 755
rect 2115 725 2290 735
rect 2115 630 2155 725
rect 1325 620 2155 630
rect 1325 600 1335 620
rect 1390 600 1820 620
rect 1875 600 2155 620
rect 1325 590 2155 600
rect -180 560 2290 570
rect -180 290 -165 560
rect -145 290 35 560
rect 55 290 235 560
rect 255 290 435 560
rect 455 290 635 560
rect 655 290 835 560
rect 855 290 885 560
rect 905 290 935 560
rect 955 290 2255 560
rect 2275 290 2290 560
rect -180 280 2290 290
rect 1025 255 2185 265
rect 1025 235 1035 255
rect 1090 235 1595 255
rect 1650 235 2120 255
rect 2175 235 2185 255
rect 1025 225 2185 235
<< labels >>
rlabel metal1 -180 1465 -180 1465 7 VP
port 1 w
rlabel metal1 -180 425 -180 425 7 VN
port 2 w
rlabel locali -180 660 -180 660 7 Vbn
port 6 w
rlabel locali -180 1305 -180 1305 7 Vbp
port 3 w
rlabel locali 2290 670 2290 670 3 Vcn
port 9 e
rlabel metal1 -180 1180 -180 1180 7 V1
port 4 w
rlabel metal1 -180 725 -180 725 7 V2
port 5 w
rlabel metal1 2290 745 2290 745 3 Vout
port 8 e
rlabel locali 2055 1690 2055 1690 3 Vcp
port 7 e
<< end >>
