magic
tech sky130A
timestamp 1616553223
<< nwell >>
rect -980 1350 -940 1450
rect -980 1205 1110 1350
rect -855 1120 -715 1205
rect 1275 1190 1480 1210
rect -970 785 -915 805
<< locali >>
rect -980 2415 -915 2425
rect -980 2395 -970 2415
rect -925 2395 -915 2415
rect -980 2385 -915 2395
rect -1060 2020 -950 2115
rect -1060 80 -1040 2020
rect -1020 1980 -975 2000
rect 985 1980 1170 2000
rect -1020 190 -1000 1980
rect 1045 1880 1130 1920
rect -980 1235 -940 1300
rect 1110 1240 1130 1880
rect 1150 1280 1170 1980
rect 1150 1260 1295 1280
rect -980 825 -960 1235
rect 1110 1220 1255 1240
rect 1215 1180 1255 1220
rect 1275 1210 1295 1260
rect 1275 1190 1480 1210
rect -980 805 -905 815
rect -980 785 -970 805
rect -915 785 -905 805
rect -980 775 -905 785
rect 1460 200 1480 1190
rect -1020 180 -940 190
rect -1020 160 -1010 180
rect -950 160 -940 180
rect 1450 160 1490 200
rect -1020 150 -940 160
rect -1060 5 -975 80
<< viali >>
rect -970 2395 -925 2415
rect -970 785 -915 805
rect -1010 160 -950 180
<< metal1 >>
rect -1060 2415 -915 2425
rect -1060 2395 -970 2415
rect -925 2395 -915 2415
rect -1060 2385 -915 2395
rect -1060 1530 -960 1820
rect -1060 1350 -915 1390
rect -855 1120 -715 1350
rect -1060 805 -905 815
rect -1060 785 -970 805
rect -915 785 -905 805
rect -1060 775 -905 785
rect -1060 670 -905 710
rect -1060 215 -905 255
rect 1470 235 1490 275
rect -1060 180 -940 190
rect -1060 160 -1010 180
rect -950 160 -940 180
rect -1060 150 -940 160
rect -1060 -210 -935 80
use fcdiffamp  fcdiffamp_0
timestamp 1616490615
transform 1 0 -800 0 1 -490
box -180 220 2290 1710
use biasgen  biasgen_0
timestamp 1616520849
transform 1 0 -1040 0 1 2735
box 60 -1500 2150 -150
<< labels >>
rlabel metal1 -1060 2405 -1060 2405 7 I1p
rlabel metal1 -1060 1675 -1060 1675 7 VP
rlabel metal1 -1060 1370 -1060 1370 7 I1n
rlabel metal1 -1060 690 -1060 690 7 V1
rlabel metal1 -1060 235 -1060 235 7 V2
rlabel metal1 -1060 -65 -1060 -65 7 VN
rlabel metal1 1490 255 1490 255 3 Vout
rlabel metal1 -1060 170 -1060 170 7 Vbn
rlabel metal1 -1060 795 -1060 795 7 Vbp
<< end >>
