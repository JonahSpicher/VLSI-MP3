magic
tech sky130A
timestamp 1616573441
<< nwell >>
rect 60 -1495 2150 -890
rect 60 -1500 165 -1495
<< nmos >>
rect 230 -260 280 -185
rect 330 -260 380 -185
rect 430 -260 480 -185
rect 530 -260 580 -185
rect 630 -260 680 -185
rect 730 -260 780 -185
rect 830 -260 880 -185
rect 930 -260 980 -185
rect 1030 -260 1080 -185
rect 1230 -260 1280 -185
rect 1330 -260 1380 -185
rect 1430 -260 1480 -185
rect 1530 -260 1580 -185
rect 1630 -260 1680 -185
rect 1730 -260 1780 -185
rect 1830 -260 1880 -185
rect 1930 -260 1980 -185
rect 2030 -260 2080 -185
rect 130 -720 180 -420
rect 230 -720 280 -420
rect 330 -720 380 -420
rect 430 -720 480 -420
rect 530 -720 580 -420
rect 630 -720 680 -420
rect 730 -720 780 -420
rect 830 -720 880 -420
rect 930 -720 980 -420
rect 1030 -720 1080 -420
rect 1130 -720 1180 -420
rect 1230 -720 1280 -420
rect 1330 -720 1380 -420
rect 1430 -720 1480 -420
rect 1530 -720 1580 -420
rect 1630 -720 1680 -420
rect 1730 -720 1780 -420
rect 1830 -720 1880 -420
rect 1930 -720 1980 -420
rect 2030 -720 2080 -420
<< pmos >>
rect 130 -1210 180 -910
rect 230 -1210 280 -910
rect 330 -1210 380 -910
rect 430 -1210 480 -910
rect 530 -1210 580 -910
rect 630 -1210 680 -910
rect 730 -1210 780 -910
rect 830 -1210 880 -910
rect 930 -1210 980 -910
rect 1030 -1210 1080 -910
rect 1130 -1210 1180 -910
rect 1230 -1210 1280 -910
rect 1330 -1210 1380 -910
rect 1430 -1210 1480 -910
rect 1530 -1210 1580 -910
rect 1630 -1210 1680 -910
rect 1730 -1210 1780 -910
rect 1830 -1210 1880 -910
rect 1930 -1210 1980 -910
rect 2030 -1210 2080 -910
rect 230 -1455 280 -1380
rect 330 -1455 380 -1380
rect 430 -1455 480 -1380
rect 530 -1455 580 -1380
rect 630 -1455 680 -1380
rect 730 -1455 780 -1380
rect 830 -1455 880 -1380
rect 930 -1455 980 -1380
rect 1030 -1455 1080 -1380
rect 1230 -1455 1280 -1380
rect 1330 -1455 1380 -1380
rect 1430 -1455 1480 -1380
rect 1530 -1455 1580 -1380
rect 1630 -1455 1680 -1380
rect 1730 -1455 1780 -1380
rect 1830 -1455 1880 -1380
rect 1930 -1455 1980 -1380
rect 2030 -1455 2080 -1380
<< ndiff >>
rect 180 -200 230 -185
rect 180 -245 195 -200
rect 215 -245 230 -200
rect 180 -260 230 -245
rect 280 -200 330 -185
rect 280 -245 295 -200
rect 315 -245 330 -200
rect 280 -260 330 -245
rect 380 -200 430 -185
rect 380 -245 395 -200
rect 415 -245 430 -200
rect 380 -260 430 -245
rect 480 -200 530 -185
rect 480 -245 495 -200
rect 515 -245 530 -200
rect 480 -260 530 -245
rect 580 -200 630 -185
rect 580 -245 595 -200
rect 615 -245 630 -200
rect 580 -260 630 -245
rect 680 -200 730 -185
rect 680 -245 695 -200
rect 715 -245 730 -200
rect 680 -260 730 -245
rect 780 -200 830 -185
rect 780 -245 795 -200
rect 815 -245 830 -200
rect 780 -260 830 -245
rect 880 -200 930 -185
rect 880 -245 895 -200
rect 915 -245 930 -200
rect 880 -260 930 -245
rect 980 -200 1030 -185
rect 980 -245 995 -200
rect 1015 -245 1030 -200
rect 980 -260 1030 -245
rect 1080 -200 1130 -185
rect 1180 -200 1230 -185
rect 1080 -245 1095 -200
rect 1115 -245 1130 -200
rect 1180 -245 1195 -200
rect 1215 -245 1230 -200
rect 1080 -260 1130 -245
rect 1180 -260 1230 -245
rect 1280 -200 1330 -185
rect 1280 -245 1295 -200
rect 1315 -245 1330 -200
rect 1280 -260 1330 -245
rect 1380 -200 1430 -185
rect 1380 -245 1395 -200
rect 1415 -245 1430 -200
rect 1380 -260 1430 -245
rect 1480 -200 1530 -185
rect 1480 -245 1495 -200
rect 1515 -245 1530 -200
rect 1480 -260 1530 -245
rect 1580 -200 1630 -185
rect 1580 -245 1595 -200
rect 1615 -245 1630 -200
rect 1580 -260 1630 -245
rect 1680 -200 1730 -185
rect 1680 -245 1695 -200
rect 1715 -245 1730 -200
rect 1680 -260 1730 -245
rect 1780 -200 1830 -185
rect 1780 -245 1795 -200
rect 1815 -245 1830 -200
rect 1780 -260 1830 -245
rect 1880 -200 1930 -185
rect 1880 -245 1895 -200
rect 1915 -245 1930 -200
rect 1880 -260 1930 -245
rect 1980 -200 2030 -185
rect 1980 -245 1995 -200
rect 2015 -245 2030 -200
rect 1980 -260 2030 -245
rect 2080 -200 2130 -185
rect 2080 -245 2095 -200
rect 2115 -245 2130 -200
rect 2080 -260 2130 -245
rect 80 -435 130 -420
rect 80 -705 95 -435
rect 115 -705 130 -435
rect 80 -720 130 -705
rect 180 -435 230 -420
rect 180 -705 195 -435
rect 215 -705 230 -435
rect 180 -720 230 -705
rect 280 -435 330 -420
rect 280 -705 295 -435
rect 315 -705 330 -435
rect 280 -720 330 -705
rect 380 -435 430 -420
rect 380 -705 395 -435
rect 415 -705 430 -435
rect 380 -720 430 -705
rect 480 -435 530 -420
rect 480 -705 495 -435
rect 515 -705 530 -435
rect 480 -720 530 -705
rect 580 -435 630 -420
rect 580 -705 595 -435
rect 615 -705 630 -435
rect 580 -720 630 -705
rect 680 -435 730 -420
rect 680 -705 695 -435
rect 715 -705 730 -435
rect 680 -720 730 -705
rect 780 -435 830 -420
rect 780 -705 795 -435
rect 815 -705 830 -435
rect 780 -720 830 -705
rect 880 -435 930 -420
rect 880 -705 895 -435
rect 915 -705 930 -435
rect 880 -720 930 -705
rect 980 -435 1030 -420
rect 980 -705 995 -435
rect 1015 -705 1030 -435
rect 980 -720 1030 -705
rect 1080 -435 1130 -420
rect 1080 -705 1095 -435
rect 1115 -705 1130 -435
rect 1080 -720 1130 -705
rect 1180 -435 1230 -420
rect 1180 -705 1195 -435
rect 1215 -705 1230 -435
rect 1180 -720 1230 -705
rect 1280 -435 1330 -420
rect 1280 -705 1295 -435
rect 1315 -705 1330 -435
rect 1280 -720 1330 -705
rect 1380 -435 1430 -420
rect 1380 -705 1395 -435
rect 1415 -705 1430 -435
rect 1380 -720 1430 -705
rect 1480 -435 1530 -420
rect 1480 -705 1495 -435
rect 1515 -705 1530 -435
rect 1480 -720 1530 -705
rect 1580 -435 1630 -420
rect 1580 -705 1595 -435
rect 1615 -705 1630 -435
rect 1580 -720 1630 -705
rect 1680 -435 1730 -420
rect 1680 -705 1695 -435
rect 1715 -705 1730 -435
rect 1680 -720 1730 -705
rect 1780 -435 1830 -420
rect 1780 -705 1795 -435
rect 1815 -705 1830 -435
rect 1780 -720 1830 -705
rect 1880 -435 1930 -420
rect 1880 -705 1895 -435
rect 1915 -705 1930 -435
rect 1880 -720 1930 -705
rect 1980 -435 2030 -420
rect 1980 -705 1995 -435
rect 2015 -705 2030 -435
rect 1980 -720 2030 -705
rect 2080 -435 2130 -420
rect 2080 -705 2095 -435
rect 2115 -705 2130 -435
rect 2080 -720 2130 -705
<< pdiff >>
rect 80 -925 130 -910
rect 80 -1195 95 -925
rect 115 -1195 130 -925
rect 80 -1210 130 -1195
rect 180 -925 230 -910
rect 180 -1195 195 -925
rect 215 -1195 230 -925
rect 180 -1210 230 -1195
rect 280 -925 330 -910
rect 280 -1195 295 -925
rect 315 -1195 330 -925
rect 280 -1210 330 -1195
rect 380 -925 430 -910
rect 380 -1195 395 -925
rect 415 -1195 430 -925
rect 380 -1210 430 -1195
rect 480 -925 530 -910
rect 480 -1195 495 -925
rect 515 -1195 530 -925
rect 480 -1210 530 -1195
rect 580 -925 630 -910
rect 580 -1195 595 -925
rect 615 -1195 630 -925
rect 580 -1210 630 -1195
rect 680 -925 730 -910
rect 680 -1195 695 -925
rect 715 -1195 730 -925
rect 680 -1210 730 -1195
rect 780 -925 830 -910
rect 780 -1195 795 -925
rect 815 -1195 830 -925
rect 780 -1210 830 -1195
rect 880 -925 930 -910
rect 880 -1195 895 -925
rect 915 -1195 930 -925
rect 880 -1210 930 -1195
rect 980 -925 1030 -910
rect 980 -1195 995 -925
rect 1015 -1195 1030 -925
rect 980 -1210 1030 -1195
rect 1080 -925 1130 -910
rect 1080 -1195 1095 -925
rect 1115 -1195 1130 -925
rect 1080 -1210 1130 -1195
rect 1180 -925 1230 -910
rect 1180 -1195 1195 -925
rect 1215 -1195 1230 -925
rect 1180 -1210 1230 -1195
rect 1280 -925 1330 -910
rect 1280 -1195 1295 -925
rect 1315 -1195 1330 -925
rect 1280 -1210 1330 -1195
rect 1380 -925 1430 -910
rect 1380 -1195 1395 -925
rect 1415 -1195 1430 -925
rect 1380 -1210 1430 -1195
rect 1480 -925 1530 -910
rect 1480 -1195 1495 -925
rect 1515 -1195 1530 -925
rect 1480 -1210 1530 -1195
rect 1580 -925 1630 -910
rect 1580 -1195 1595 -925
rect 1615 -1195 1630 -925
rect 1580 -1210 1630 -1195
rect 1680 -925 1730 -910
rect 1680 -1195 1695 -925
rect 1715 -1195 1730 -925
rect 1680 -1210 1730 -1195
rect 1780 -925 1830 -910
rect 1780 -1195 1795 -925
rect 1815 -1195 1830 -925
rect 1780 -1210 1830 -1195
rect 1880 -925 1930 -910
rect 1880 -1195 1895 -925
rect 1915 -1195 1930 -925
rect 1880 -1210 1930 -1195
rect 1980 -925 2030 -910
rect 1980 -1195 1995 -925
rect 2015 -1195 2030 -925
rect 1980 -1210 2030 -1195
rect 2080 -925 2130 -910
rect 2080 -1195 2095 -925
rect 2115 -1195 2130 -925
rect 2080 -1210 2130 -1195
rect 180 -1395 230 -1380
rect 180 -1440 195 -1395
rect 215 -1440 230 -1395
rect 180 -1455 230 -1440
rect 280 -1395 330 -1380
rect 280 -1440 295 -1395
rect 315 -1440 330 -1395
rect 280 -1455 330 -1440
rect 380 -1395 430 -1380
rect 380 -1440 395 -1395
rect 415 -1440 430 -1395
rect 380 -1455 430 -1440
rect 480 -1395 530 -1380
rect 480 -1440 495 -1395
rect 515 -1440 530 -1395
rect 480 -1455 530 -1440
rect 580 -1395 630 -1380
rect 580 -1440 595 -1395
rect 615 -1440 630 -1395
rect 580 -1455 630 -1440
rect 680 -1395 730 -1380
rect 680 -1440 695 -1395
rect 715 -1440 730 -1395
rect 680 -1455 730 -1440
rect 780 -1395 830 -1380
rect 780 -1440 795 -1395
rect 815 -1440 830 -1395
rect 780 -1455 830 -1440
rect 880 -1395 930 -1380
rect 880 -1440 895 -1395
rect 915 -1440 930 -1395
rect 880 -1455 930 -1440
rect 980 -1395 1030 -1380
rect 980 -1440 995 -1395
rect 1015 -1440 1030 -1395
rect 980 -1455 1030 -1440
rect 1080 -1395 1130 -1380
rect 1180 -1395 1230 -1380
rect 1080 -1440 1095 -1395
rect 1115 -1440 1130 -1395
rect 1180 -1440 1195 -1395
rect 1215 -1440 1230 -1395
rect 1080 -1455 1130 -1440
rect 1180 -1455 1230 -1440
rect 1280 -1395 1330 -1380
rect 1280 -1440 1295 -1395
rect 1315 -1440 1330 -1395
rect 1280 -1455 1330 -1440
rect 1380 -1395 1430 -1380
rect 1380 -1440 1395 -1395
rect 1415 -1440 1430 -1395
rect 1380 -1455 1430 -1440
rect 1480 -1395 1530 -1380
rect 1480 -1440 1495 -1395
rect 1515 -1440 1530 -1395
rect 1480 -1455 1530 -1440
rect 1580 -1395 1630 -1380
rect 1580 -1440 1595 -1395
rect 1615 -1440 1630 -1395
rect 1580 -1455 1630 -1440
rect 1680 -1395 1730 -1380
rect 1680 -1440 1695 -1395
rect 1715 -1440 1730 -1395
rect 1680 -1455 1730 -1440
rect 1780 -1395 1830 -1380
rect 1780 -1440 1795 -1395
rect 1815 -1440 1830 -1395
rect 1780 -1455 1830 -1440
rect 1880 -1395 1930 -1380
rect 1880 -1440 1895 -1395
rect 1915 -1440 1930 -1395
rect 1880 -1455 1930 -1440
rect 1980 -1395 2030 -1380
rect 1980 -1440 1995 -1395
rect 2015 -1440 2030 -1395
rect 1980 -1455 2030 -1440
rect 2080 -1395 2130 -1380
rect 2080 -1440 2095 -1395
rect 2115 -1440 2130 -1395
rect 2080 -1455 2130 -1440
<< ndiffc >>
rect 195 -245 215 -200
rect 295 -245 315 -200
rect 395 -245 415 -200
rect 495 -245 515 -200
rect 595 -245 615 -200
rect 695 -245 715 -200
rect 795 -245 815 -200
rect 895 -245 915 -200
rect 995 -245 1015 -200
rect 1095 -245 1115 -200
rect 1195 -245 1215 -200
rect 1295 -245 1315 -200
rect 1395 -245 1415 -200
rect 1495 -245 1515 -200
rect 1595 -245 1615 -200
rect 1695 -245 1715 -200
rect 1795 -245 1815 -200
rect 1895 -245 1915 -200
rect 1995 -245 2015 -200
rect 2095 -245 2115 -200
rect 95 -705 115 -435
rect 195 -705 215 -435
rect 295 -705 315 -435
rect 395 -705 415 -435
rect 495 -705 515 -435
rect 595 -705 615 -435
rect 695 -705 715 -435
rect 795 -705 815 -435
rect 895 -705 915 -435
rect 995 -705 1015 -435
rect 1095 -705 1115 -435
rect 1195 -705 1215 -435
rect 1295 -705 1315 -435
rect 1395 -705 1415 -435
rect 1495 -705 1515 -435
rect 1595 -705 1615 -435
rect 1695 -705 1715 -435
rect 1795 -705 1815 -435
rect 1895 -705 1915 -435
rect 1995 -705 2015 -435
rect 2095 -705 2115 -435
<< pdiffc >>
rect 95 -1195 115 -925
rect 195 -1195 215 -925
rect 295 -1195 315 -925
rect 395 -1195 415 -925
rect 495 -1195 515 -925
rect 595 -1195 615 -925
rect 695 -1195 715 -925
rect 795 -1195 815 -925
rect 895 -1195 915 -925
rect 995 -1195 1015 -925
rect 1095 -1195 1115 -925
rect 1195 -1195 1215 -925
rect 1295 -1195 1315 -925
rect 1395 -1195 1415 -925
rect 1495 -1195 1515 -925
rect 1595 -1195 1615 -925
rect 1695 -1195 1715 -925
rect 1795 -1195 1815 -925
rect 1895 -1195 1915 -925
rect 1995 -1195 2015 -925
rect 2095 -1195 2115 -925
rect 195 -1440 215 -1395
rect 295 -1440 315 -1395
rect 395 -1440 415 -1395
rect 495 -1440 515 -1395
rect 595 -1440 615 -1395
rect 695 -1440 715 -1395
rect 795 -1440 815 -1395
rect 895 -1440 915 -1395
rect 995 -1440 1015 -1395
rect 1095 -1440 1115 -1395
rect 1195 -1440 1215 -1395
rect 1295 -1440 1315 -1395
rect 1395 -1440 1415 -1395
rect 1495 -1440 1515 -1395
rect 1595 -1440 1615 -1395
rect 1695 -1440 1715 -1395
rect 1795 -1440 1815 -1395
rect 1895 -1440 1915 -1395
rect 1995 -1440 2015 -1395
rect 2095 -1440 2115 -1395
<< psubdiff >>
rect 1130 -200 1180 -185
rect 1130 -245 1145 -200
rect 1165 -245 1180 -200
rect 1130 -260 1180 -245
<< nsubdiff >>
rect 1130 -1395 1180 -1380
rect 1130 -1440 1145 -1395
rect 1165 -1440 1180 -1395
rect 1130 -1455 1180 -1440
<< psubdiffcont >>
rect 1145 -245 1165 -200
<< nsubdiffcont >>
rect 1145 -1440 1165 -1395
<< poly >>
rect 230 -185 280 -170
rect 330 -185 380 -170
rect 430 -185 480 -170
rect 530 -185 580 -170
rect 630 -185 680 -170
rect 730 -185 780 -170
rect 830 -185 880 -170
rect 930 -185 980 -170
rect 1030 -185 1080 -170
rect 1230 -185 1280 -170
rect 1330 -185 1380 -170
rect 1430 -185 1480 -170
rect 1530 -185 1580 -170
rect 1630 -185 1680 -170
rect 1730 -185 1780 -170
rect 1830 -185 1880 -170
rect 1930 -185 1980 -170
rect 2030 -185 2080 -170
rect 230 -275 280 -260
rect 330 -270 380 -260
rect 430 -270 480 -260
rect 530 -270 580 -260
rect 630 -270 680 -260
rect 730 -270 780 -260
rect 830 -270 880 -260
rect 930 -270 980 -260
rect 1030 -270 1080 -260
rect 1230 -270 1280 -260
rect 1330 -270 1380 -260
rect 1430 -270 1480 -260
rect 1530 -270 1580 -260
rect 1630 -270 1680 -260
rect 1730 -270 1780 -260
rect 1830 -270 1880 -260
rect 1930 -270 1980 -260
rect 230 -280 270 -275
rect 230 -300 240 -280
rect 260 -300 270 -280
rect 330 -285 1980 -270
rect 2030 -275 2080 -260
rect 2040 -280 2080 -275
rect 230 -310 270 -300
rect 1230 -305 1240 -285
rect 1260 -305 1270 -285
rect 1230 -315 1270 -305
rect 2040 -300 2050 -280
rect 2070 -300 2080 -280
rect 2040 -310 2080 -300
rect 130 -380 170 -370
rect 130 -400 140 -380
rect 160 -400 170 -380
rect 130 -405 170 -400
rect 230 -380 270 -370
rect 230 -400 240 -380
rect 260 -395 270 -380
rect 585 -380 625 -370
rect 585 -395 595 -380
rect 260 -400 595 -395
rect 615 -395 625 -380
rect 940 -380 980 -370
rect 940 -395 950 -380
rect 615 -400 950 -395
rect 970 -400 980 -380
rect 1085 -380 1125 -370
rect 1085 -395 1095 -380
rect 130 -420 180 -405
rect 230 -410 980 -400
rect 230 -420 280 -410
rect 330 -420 380 -410
rect 430 -420 480 -410
rect 530 -420 580 -410
rect 630 -420 680 -410
rect 730 -420 780 -410
rect 830 -420 880 -410
rect 930 -420 980 -410
rect 1030 -400 1095 -395
rect 1115 -395 1125 -380
rect 1230 -380 1270 -370
rect 1115 -400 1180 -395
rect 1030 -410 1180 -400
rect 1030 -420 1080 -410
rect 1130 -420 1180 -410
rect 1230 -400 1240 -380
rect 1260 -400 1270 -380
rect 1585 -380 1625 -370
rect 1585 -395 1595 -380
rect 1230 -405 1270 -400
rect 1530 -400 1595 -395
rect 1615 -395 1625 -380
rect 1940 -380 1980 -370
rect 1615 -400 1680 -395
rect 1230 -420 1280 -405
rect 1330 -420 1380 -405
rect 1430 -420 1480 -405
rect 1530 -410 1680 -400
rect 1940 -400 1950 -380
rect 1970 -400 1980 -380
rect 1940 -405 1980 -400
rect 2040 -380 2080 -370
rect 2040 -400 2050 -380
rect 2070 -400 2080 -380
rect 2040 -405 2080 -400
rect 1530 -420 1580 -410
rect 1630 -420 1680 -410
rect 1730 -420 1780 -405
rect 1830 -420 1880 -405
rect 1930 -420 1980 -405
rect 2030 -420 2080 -405
rect 130 -735 180 -720
rect 230 -735 280 -720
rect 330 -735 380 -720
rect 430 -735 480 -720
rect 530 -735 580 -720
rect 630 -735 680 -720
rect 730 -735 780 -720
rect 830 -735 880 -720
rect 930 -735 980 -720
rect 1030 -735 1080 -720
rect 1130 -735 1180 -720
rect 1230 -735 1280 -720
rect 1330 -730 1380 -720
rect 1430 -730 1480 -720
rect 1330 -740 1480 -730
rect 1530 -735 1580 -720
rect 1630 -735 1680 -720
rect 1730 -730 1780 -720
rect 1830 -730 1880 -720
rect 1330 -745 1395 -740
rect 1385 -760 1395 -745
rect 1415 -760 1480 -740
rect 1730 -740 1880 -730
rect 1930 -735 1980 -720
rect 2030 -735 2080 -720
rect 1730 -760 1795 -740
rect 1815 -750 1880 -740
rect 1815 -760 1825 -750
rect 1385 -775 1825 -760
rect 1810 -830 1825 -775
rect 1785 -840 1825 -830
rect 240 -865 970 -855
rect 240 -885 250 -865
rect 270 -870 595 -865
rect 270 -885 280 -870
rect 240 -895 280 -885
rect 530 -885 595 -870
rect 615 -870 940 -865
rect 615 -885 680 -870
rect 130 -910 180 -895
rect 230 -910 280 -895
rect 330 -910 380 -895
rect 430 -910 480 -895
rect 530 -900 680 -885
rect 930 -885 940 -870
rect 960 -885 970 -865
rect 1785 -860 1795 -840
rect 1815 -860 1825 -840
rect 1785 -870 1825 -860
rect 930 -895 970 -885
rect 530 -910 580 -900
rect 630 -910 680 -900
rect 730 -910 780 -895
rect 830 -910 880 -895
rect 930 -910 980 -895
rect 1030 -910 1080 -895
rect 1130 -910 1180 -895
rect 1230 -910 1280 -895
rect 1330 -910 1380 -895
rect 1430 -910 1480 -895
rect 1530 -910 1580 -895
rect 1630 -910 1680 -895
rect 1730 -910 1780 -895
rect 1830 -910 1880 -895
rect 1930 -910 1980 -895
rect 2030 -910 2080 -895
rect 130 -1225 180 -1210
rect 230 -1225 280 -1210
rect 330 -1220 380 -1210
rect 430 -1220 480 -1210
rect 130 -1235 170 -1225
rect 330 -1235 480 -1220
rect 530 -1225 580 -1210
rect 630 -1225 680 -1210
rect 730 -1220 780 -1210
rect 830 -1220 880 -1210
rect 130 -1255 140 -1235
rect 160 -1250 170 -1235
rect 160 -1255 245 -1250
rect 130 -1265 245 -1255
rect 385 -1255 395 -1235
rect 415 -1250 480 -1235
rect 730 -1235 880 -1220
rect 930 -1225 980 -1210
rect 1030 -1220 1080 -1210
rect 1130 -1220 1180 -1210
rect 1030 -1225 1180 -1220
rect 1230 -1220 1280 -1210
rect 1330 -1220 1380 -1210
rect 1430 -1220 1480 -1210
rect 1530 -1220 1580 -1210
rect 1630 -1220 1680 -1210
rect 1730 -1220 1780 -1210
rect 1830 -1220 1880 -1210
rect 1930 -1220 1980 -1210
rect 1030 -1235 1170 -1225
rect 730 -1250 795 -1235
rect 415 -1255 795 -1250
rect 815 -1255 825 -1235
rect 1030 -1240 1140 -1235
rect 385 -1265 825 -1255
rect 1130 -1255 1140 -1240
rect 1160 -1255 1170 -1235
rect 1130 -1265 1170 -1255
rect 1230 -1235 1980 -1220
rect 2030 -1225 2080 -1210
rect 1230 -1255 1240 -1235
rect 1260 -1255 1270 -1235
rect 1230 -1265 1270 -1255
rect 1585 -1255 1595 -1235
rect 1615 -1255 1625 -1235
rect 1585 -1265 1625 -1255
rect 1940 -1255 1950 -1235
rect 1970 -1255 1980 -1235
rect 1940 -1265 1980 -1255
rect 2040 -1235 2080 -1225
rect 2040 -1255 2050 -1235
rect 2070 -1255 2080 -1235
rect 2040 -1265 2080 -1255
rect 230 -1365 245 -1265
rect 785 -1335 825 -1325
rect 785 -1355 795 -1335
rect 815 -1355 825 -1335
rect 230 -1380 280 -1365
rect 330 -1370 1980 -1355
rect 2060 -1365 2080 -1265
rect 330 -1380 380 -1370
rect 430 -1380 480 -1370
rect 530 -1380 580 -1370
rect 630 -1380 680 -1370
rect 730 -1380 780 -1370
rect 830 -1380 880 -1370
rect 930 -1380 980 -1370
rect 1030 -1380 1080 -1370
rect 1230 -1380 1280 -1370
rect 1330 -1380 1380 -1370
rect 1430 -1380 1480 -1370
rect 1530 -1380 1580 -1370
rect 1630 -1380 1680 -1370
rect 1730 -1380 1780 -1370
rect 1830 -1380 1880 -1370
rect 1930 -1380 1980 -1370
rect 2030 -1380 2080 -1365
rect 230 -1470 280 -1455
rect 330 -1470 380 -1455
rect 430 -1470 480 -1455
rect 530 -1470 580 -1455
rect 630 -1470 680 -1455
rect 730 -1470 780 -1455
rect 830 -1470 880 -1455
rect 930 -1470 980 -1455
rect 1030 -1470 1080 -1455
rect 1230 -1470 1280 -1455
rect 1330 -1470 1380 -1455
rect 1430 -1470 1480 -1455
rect 1530 -1470 1580 -1455
rect 1630 -1470 1680 -1455
rect 1730 -1470 1780 -1455
rect 1830 -1470 1880 -1455
rect 1930 -1470 1980 -1455
rect 2030 -1470 2080 -1455
<< polycont >>
rect 240 -300 260 -280
rect 1240 -305 1260 -285
rect 2050 -300 2070 -280
rect 140 -400 160 -380
rect 240 -400 260 -380
rect 595 -400 615 -380
rect 950 -400 970 -380
rect 1095 -400 1115 -380
rect 1240 -400 1260 -380
rect 1595 -400 1615 -380
rect 1950 -400 1970 -380
rect 2050 -400 2070 -380
rect 1395 -760 1415 -740
rect 1795 -760 1815 -740
rect 250 -885 270 -865
rect 595 -885 615 -865
rect 940 -885 960 -865
rect 1795 -860 1815 -840
rect 140 -1255 160 -1235
rect 395 -1255 415 -1235
rect 795 -1255 815 -1235
rect 1140 -1255 1160 -1235
rect 1240 -1255 1260 -1235
rect 1595 -1255 1615 -1235
rect 1950 -1255 1970 -1235
rect 2050 -1255 2070 -1235
rect 795 -1355 815 -1335
<< locali >>
rect 405 -170 1905 -150
rect 405 -190 425 -170
rect 605 -190 625 -170
rect 805 -190 825 -170
rect 1005 -190 1025 -170
rect 1285 -190 1305 -170
rect 1485 -190 1505 -170
rect 1685 -190 1705 -170
rect 1885 -190 1905 -170
rect 185 -200 225 -190
rect 185 -245 195 -200
rect 215 -245 225 -200
rect 185 -255 225 -245
rect 285 -200 325 -190
rect 285 -245 295 -200
rect 315 -245 325 -200
rect 285 -255 325 -245
rect 385 -200 425 -190
rect 385 -245 395 -200
rect 415 -245 425 -200
rect 385 -255 425 -245
rect 485 -200 525 -190
rect 485 -245 495 -200
rect 515 -245 525 -200
rect 485 -255 525 -245
rect 585 -200 625 -190
rect 585 -245 595 -200
rect 615 -245 625 -200
rect 585 -255 625 -245
rect 685 -200 725 -190
rect 685 -245 695 -200
rect 715 -245 725 -200
rect 685 -255 725 -245
rect 785 -200 825 -190
rect 785 -245 795 -200
rect 815 -245 825 -200
rect 785 -255 825 -245
rect 885 -200 925 -190
rect 885 -245 895 -200
rect 915 -245 925 -200
rect 885 -255 925 -245
rect 985 -200 1025 -190
rect 985 -245 995 -200
rect 1015 -245 1025 -200
rect 985 -255 1025 -245
rect 1085 -200 1225 -190
rect 1085 -245 1095 -200
rect 1115 -245 1145 -200
rect 1165 -245 1195 -200
rect 1215 -245 1225 -200
rect 1085 -255 1225 -245
rect 1285 -200 1325 -190
rect 1285 -245 1295 -200
rect 1315 -245 1325 -200
rect 1285 -255 1325 -245
rect 1385 -200 1425 -190
rect 1385 -245 1395 -200
rect 1415 -245 1425 -200
rect 1385 -255 1425 -245
rect 1485 -200 1525 -190
rect 1485 -245 1495 -200
rect 1515 -245 1525 -200
rect 1485 -255 1525 -245
rect 1585 -200 1625 -190
rect 1585 -245 1595 -200
rect 1615 -245 1625 -200
rect 1585 -255 1625 -245
rect 1685 -200 1725 -190
rect 1685 -245 1695 -200
rect 1715 -245 1725 -200
rect 1685 -255 1725 -245
rect 1785 -200 1825 -190
rect 1785 -245 1795 -200
rect 1815 -245 1825 -200
rect 1785 -255 1825 -245
rect 1885 -200 1925 -190
rect 1885 -245 1895 -200
rect 1915 -245 1925 -200
rect 1885 -255 1925 -245
rect 1985 -200 2025 -190
rect 1985 -245 1995 -200
rect 2015 -245 2025 -200
rect 1985 -255 2025 -245
rect 2085 -200 2125 -190
rect 2085 -245 2095 -200
rect 2115 -245 2125 -200
rect 2085 -255 2125 -245
rect 205 -270 225 -255
rect 205 -280 270 -270
rect 205 -290 240 -280
rect 230 -300 240 -290
rect 260 -300 270 -280
rect 230 -310 270 -300
rect 1230 -285 1270 -275
rect 1230 -305 1240 -285
rect 1260 -305 1270 -285
rect 1230 -315 1270 -305
rect 1230 -330 1250 -315
rect 60 -350 1250 -330
rect 1230 -370 1250 -350
rect 1305 -330 1325 -255
rect 2085 -270 2105 -255
rect 2040 -280 2105 -270
rect 2040 -300 2050 -280
rect 2070 -290 2105 -280
rect 2070 -300 2080 -290
rect 2040 -310 2080 -300
rect 1305 -350 1905 -330
rect 130 -380 170 -370
rect 130 -390 140 -380
rect 105 -400 140 -390
rect 160 -400 170 -380
rect 230 -380 270 -370
rect 230 -390 240 -380
rect 105 -410 170 -400
rect 205 -400 240 -390
rect 260 -400 270 -380
rect 205 -410 270 -400
rect 585 -380 625 -370
rect 585 -400 595 -380
rect 615 -400 625 -380
rect 105 -425 125 -410
rect 205 -425 225 -410
rect 85 -435 125 -425
rect 85 -705 95 -435
rect 115 -705 125 -435
rect 85 -715 125 -705
rect 185 -435 225 -425
rect 185 -705 195 -435
rect 215 -705 225 -435
rect 185 -715 225 -705
rect 285 -435 325 -425
rect 285 -705 295 -435
rect 315 -705 325 -435
rect 285 -715 325 -705
rect 385 -435 425 -425
rect 385 -705 395 -435
rect 415 -705 425 -435
rect 385 -715 425 -705
rect 485 -435 525 -425
rect 485 -705 495 -435
rect 515 -705 525 -435
rect 485 -715 525 -705
rect 585 -435 625 -400
rect 940 -380 980 -370
rect 940 -400 950 -380
rect 970 -390 980 -380
rect 1085 -380 1125 -370
rect 970 -400 1005 -390
rect 940 -410 1005 -400
rect 985 -425 1005 -410
rect 1085 -400 1095 -380
rect 1115 -400 1125 -380
rect 1230 -380 1270 -370
rect 1230 -390 1240 -380
rect 585 -705 595 -435
rect 615 -705 625 -435
rect 585 -715 625 -705
rect 685 -435 725 -425
rect 685 -705 695 -435
rect 715 -705 725 -435
rect 685 -715 725 -705
rect 785 -435 825 -425
rect 785 -705 795 -435
rect 815 -705 825 -435
rect 785 -715 825 -705
rect 885 -435 925 -425
rect 885 -705 895 -435
rect 915 -705 925 -435
rect 885 -715 925 -705
rect 985 -435 1025 -425
rect 985 -705 995 -435
rect 1015 -705 1025 -435
rect 985 -715 1025 -705
rect 1085 -435 1125 -400
rect 1205 -400 1240 -390
rect 1260 -400 1270 -380
rect 1205 -410 1270 -400
rect 1205 -425 1225 -410
rect 1305 -425 1325 -350
rect 1485 -425 1505 -350
rect 1585 -380 1625 -370
rect 1585 -400 1595 -380
rect 1615 -400 1625 -380
rect 1085 -705 1095 -435
rect 1115 -705 1125 -435
rect 1085 -715 1125 -705
rect 1185 -435 1225 -425
rect 1185 -705 1195 -435
rect 1215 -705 1225 -435
rect 1185 -715 1225 -705
rect 1285 -435 1325 -425
rect 1285 -705 1295 -435
rect 1315 -705 1325 -435
rect 1285 -715 1325 -705
rect 1385 -435 1425 -425
rect 1385 -705 1395 -435
rect 1415 -705 1425 -435
rect 185 -735 205 -715
rect 405 -735 425 -715
rect 785 -735 805 -715
rect 60 -755 205 -735
rect 260 -755 805 -735
rect 260 -855 280 -755
rect 1205 -790 1225 -715
rect 1385 -740 1425 -705
rect 1485 -435 1525 -425
rect 1485 -705 1495 -435
rect 1515 -705 1525 -435
rect 1485 -715 1525 -705
rect 1585 -435 1625 -400
rect 1585 -705 1595 -435
rect 1615 -705 1625 -435
rect 1585 -715 1625 -705
rect 1685 -425 1705 -350
rect 1885 -425 1905 -350
rect 1940 -380 1980 -370
rect 1940 -400 1950 -380
rect 1970 -390 1980 -380
rect 2040 -380 2080 -370
rect 1970 -400 2005 -390
rect 1940 -410 2005 -400
rect 2040 -400 2050 -380
rect 2070 -390 2080 -380
rect 2070 -400 2105 -390
rect 2040 -410 2105 -400
rect 1985 -425 2005 -410
rect 2085 -425 2105 -410
rect 1685 -435 1725 -425
rect 1685 -705 1695 -435
rect 1715 -705 1725 -435
rect 1685 -715 1725 -705
rect 1785 -435 1825 -425
rect 1785 -705 1795 -435
rect 1815 -705 1825 -435
rect 1385 -760 1395 -740
rect 1415 -760 1425 -740
rect 1385 -770 1425 -760
rect 1585 -790 1605 -715
rect 1785 -740 1825 -705
rect 1885 -435 1925 -425
rect 1885 -705 1895 -435
rect 1915 -705 1925 -435
rect 1885 -715 1925 -705
rect 1985 -435 2025 -425
rect 1985 -705 1995 -435
rect 2015 -705 2025 -435
rect 1985 -715 2025 -705
rect 2085 -435 2125 -425
rect 2085 -705 2095 -435
rect 2115 -705 2125 -435
rect 2085 -715 2125 -705
rect 1785 -760 1795 -740
rect 1815 -760 1825 -740
rect 1785 -770 1825 -760
rect 1985 -790 2005 -715
rect 1205 -810 2005 -790
rect 2025 -755 2150 -735
rect 240 -865 280 -855
rect 240 -875 250 -865
rect 205 -885 250 -875
rect 270 -885 280 -865
rect 205 -895 280 -885
rect 305 -835 905 -815
rect 2025 -830 2045 -755
rect 205 -915 225 -895
rect 305 -915 325 -835
rect 505 -915 525 -835
rect 85 -925 125 -915
rect 85 -1195 95 -925
rect 115 -1195 125 -925
rect 85 -1205 125 -1195
rect 185 -925 225 -915
rect 185 -1195 195 -925
rect 215 -1195 225 -925
rect 185 -1205 225 -1195
rect 285 -925 325 -915
rect 285 -1195 295 -925
rect 315 -1195 325 -925
rect 285 -1205 325 -1195
rect 385 -925 425 -915
rect 385 -1195 395 -925
rect 415 -1195 425 -925
rect 105 -1225 125 -1205
rect 105 -1235 170 -1225
rect 105 -1245 140 -1235
rect 130 -1255 140 -1245
rect 160 -1255 170 -1235
rect 130 -1265 170 -1255
rect 385 -1235 425 -1195
rect 485 -925 525 -915
rect 485 -1195 495 -925
rect 515 -1195 525 -925
rect 485 -1205 525 -1195
rect 585 -865 625 -855
rect 585 -885 595 -865
rect 615 -885 625 -865
rect 585 -925 625 -885
rect 585 -1195 595 -925
rect 615 -1195 625 -925
rect 585 -1205 625 -1195
rect 685 -915 705 -835
rect 885 -915 905 -835
rect 930 -840 970 -830
rect 930 -885 940 -840
rect 960 -875 970 -840
rect 1785 -840 2045 -830
rect 1785 -860 1795 -840
rect 1815 -850 2045 -840
rect 2085 -825 2150 -815
rect 2085 -845 2095 -825
rect 2140 -845 2150 -825
rect 1815 -860 1825 -850
rect 2085 -855 2150 -845
rect 1785 -870 1825 -860
rect 1785 -875 1805 -870
rect 960 -885 1005 -875
rect 930 -895 1005 -885
rect 985 -915 1005 -895
rect 1405 -895 1805 -875
rect 1405 -915 1425 -895
rect 1785 -915 1805 -895
rect 685 -925 725 -915
rect 685 -1195 695 -925
rect 715 -1195 725 -925
rect 685 -1205 725 -1195
rect 385 -1255 395 -1235
rect 415 -1255 425 -1235
rect 385 -1265 425 -1255
rect 385 -1345 405 -1265
rect 705 -1345 725 -1205
rect 785 -925 825 -915
rect 785 -1195 795 -925
rect 815 -1195 825 -925
rect 785 -1235 825 -1195
rect 885 -925 925 -915
rect 885 -1195 895 -925
rect 915 -1195 925 -925
rect 885 -1205 925 -1195
rect 985 -925 1025 -915
rect 985 -1195 995 -925
rect 1015 -1195 1025 -925
rect 985 -1205 1025 -1195
rect 1085 -925 1125 -915
rect 1085 -1195 1095 -925
rect 1115 -1195 1125 -925
rect 1085 -1205 1125 -1195
rect 1185 -925 1225 -915
rect 1185 -1195 1195 -925
rect 1215 -1195 1225 -925
rect 1185 -1205 1225 -1195
rect 1285 -925 1325 -915
rect 1285 -1195 1295 -925
rect 1315 -1195 1325 -925
rect 1285 -1205 1325 -1195
rect 1385 -925 1425 -915
rect 1385 -1195 1395 -925
rect 1415 -1195 1425 -925
rect 1385 -1205 1425 -1195
rect 1485 -925 1525 -915
rect 1485 -1195 1495 -925
rect 1515 -1195 1525 -925
rect 1485 -1205 1525 -1195
rect 1585 -925 1625 -915
rect 1585 -1195 1595 -925
rect 1615 -1195 1625 -925
rect 785 -1255 795 -1235
rect 815 -1255 825 -1235
rect 1105 -1225 1125 -1205
rect 1205 -1225 1225 -1205
rect 1105 -1235 1170 -1225
rect 1105 -1245 1140 -1235
rect 785 -1265 825 -1255
rect 1130 -1255 1140 -1245
rect 1160 -1255 1170 -1235
rect 1205 -1235 1270 -1225
rect 1205 -1245 1240 -1235
rect 1130 -1265 1170 -1255
rect 1230 -1255 1240 -1245
rect 1260 -1255 1270 -1235
rect 1230 -1265 1270 -1255
rect 1585 -1235 1625 -1195
rect 1685 -925 1725 -915
rect 1685 -1195 1695 -925
rect 1715 -1195 1725 -925
rect 1685 -1205 1725 -1195
rect 1785 -925 1825 -915
rect 1785 -1195 1795 -925
rect 1815 -1195 1825 -925
rect 1785 -1205 1825 -1195
rect 1885 -925 1925 -915
rect 1885 -1195 1895 -925
rect 1915 -1195 1925 -925
rect 1885 -1205 1925 -1195
rect 1985 -925 2025 -915
rect 1985 -1195 1995 -925
rect 2015 -1195 2025 -925
rect 1985 -1205 2025 -1195
rect 2085 -925 2125 -915
rect 2085 -1195 2095 -925
rect 2115 -1195 2125 -925
rect 2085 -1205 2125 -1195
rect 1985 -1225 2005 -1205
rect 2085 -1225 2105 -1205
rect 1585 -1255 1595 -1235
rect 1615 -1255 1625 -1235
rect 1585 -1265 1625 -1255
rect 1940 -1235 2005 -1225
rect 1940 -1255 1950 -1235
rect 1970 -1245 2005 -1235
rect 2040 -1235 2105 -1225
rect 1970 -1255 1980 -1245
rect 1940 -1265 1980 -1255
rect 2040 -1255 2050 -1235
rect 2070 -1245 2105 -1235
rect 2070 -1255 2080 -1245
rect 2040 -1265 2080 -1255
rect 805 -1325 825 -1265
rect 1230 -1285 1250 -1265
rect 1185 -1295 1250 -1285
rect 1185 -1315 1195 -1295
rect 1240 -1315 1250 -1295
rect 1185 -1325 1250 -1315
rect 60 -1355 405 -1345
rect 60 -1375 70 -1355
rect 115 -1365 405 -1355
rect 605 -1365 725 -1345
rect 785 -1335 825 -1325
rect 785 -1355 795 -1335
rect 815 -1355 825 -1335
rect 785 -1365 825 -1355
rect 115 -1375 125 -1365
rect 60 -1385 125 -1375
rect 605 -1385 625 -1365
rect 185 -1395 225 -1385
rect 60 -1445 100 -1435
rect 60 -1490 70 -1445
rect 90 -1490 100 -1445
rect 185 -1440 195 -1395
rect 215 -1440 225 -1395
rect 185 -1450 225 -1440
rect 285 -1395 325 -1385
rect 285 -1440 295 -1395
rect 315 -1440 325 -1395
rect 285 -1450 325 -1440
rect 385 -1395 425 -1385
rect 385 -1440 395 -1395
rect 415 -1440 425 -1395
rect 385 -1450 425 -1440
rect 485 -1395 525 -1385
rect 485 -1440 495 -1395
rect 515 -1440 525 -1395
rect 485 -1450 525 -1440
rect 585 -1395 625 -1385
rect 585 -1440 595 -1395
rect 615 -1440 625 -1395
rect 585 -1450 625 -1440
rect 685 -1395 725 -1385
rect 685 -1440 695 -1395
rect 715 -1440 725 -1395
rect 685 -1450 725 -1440
rect 785 -1395 825 -1385
rect 785 -1440 795 -1395
rect 815 -1440 825 -1395
rect 785 -1450 825 -1440
rect 885 -1395 925 -1385
rect 885 -1440 895 -1395
rect 915 -1440 925 -1395
rect 885 -1450 925 -1440
rect 985 -1395 1025 -1385
rect 985 -1440 995 -1395
rect 1015 -1440 1025 -1395
rect 985 -1450 1025 -1440
rect 1085 -1395 1225 -1385
rect 1085 -1440 1095 -1395
rect 1115 -1440 1145 -1395
rect 1165 -1440 1195 -1395
rect 1215 -1440 1225 -1395
rect 1085 -1450 1225 -1440
rect 1285 -1395 1325 -1385
rect 1285 -1440 1295 -1395
rect 1315 -1440 1325 -1395
rect 1285 -1450 1325 -1440
rect 1385 -1395 1425 -1385
rect 1385 -1440 1395 -1395
rect 1415 -1440 1425 -1395
rect 1385 -1450 1425 -1440
rect 1485 -1395 1525 -1385
rect 1485 -1440 1495 -1395
rect 1515 -1440 1525 -1395
rect 1485 -1450 1525 -1440
rect 1585 -1395 1625 -1385
rect 1585 -1440 1595 -1395
rect 1615 -1440 1625 -1395
rect 1585 -1450 1625 -1440
rect 1685 -1395 1725 -1385
rect 1685 -1440 1695 -1395
rect 1715 -1440 1725 -1395
rect 1685 -1450 1725 -1440
rect 1785 -1395 1825 -1385
rect 1785 -1440 1795 -1395
rect 1815 -1440 1825 -1395
rect 1785 -1450 1825 -1440
rect 1885 -1395 1925 -1385
rect 1885 -1440 1895 -1395
rect 1915 -1440 1925 -1395
rect 1885 -1450 1925 -1440
rect 1985 -1395 2025 -1385
rect 1985 -1440 1995 -1395
rect 2015 -1440 2025 -1395
rect 1985 -1450 2025 -1440
rect 2085 -1395 2125 -1385
rect 2085 -1440 2095 -1395
rect 2115 -1440 2125 -1395
rect 2085 -1450 2125 -1440
rect 405 -1470 425 -1450
rect 605 -1470 625 -1450
rect 805 -1470 825 -1450
rect 1005 -1470 1025 -1450
rect 1285 -1470 1305 -1450
rect 1485 -1470 1505 -1450
rect 1685 -1470 1705 -1450
rect 1885 -1470 1905 -1450
rect 405 -1490 1905 -1470
rect 60 -1500 100 -1490
<< viali >>
rect 195 -245 215 -200
rect 295 -245 315 -200
rect 495 -245 515 -200
rect 695 -245 715 -200
rect 895 -245 915 -200
rect 1095 -245 1115 -200
rect 1145 -245 1165 -200
rect 1195 -245 1215 -200
rect 1395 -245 1415 -200
rect 1595 -245 1615 -200
rect 1795 -245 1815 -200
rect 1995 -245 2015 -200
rect 2095 -245 2115 -200
rect 95 -705 115 -435
rect 295 -705 315 -435
rect 495 -705 515 -435
rect 695 -705 715 -435
rect 895 -705 915 -435
rect 1095 -705 1115 -435
rect 2095 -705 2115 -435
rect 95 -1195 115 -925
rect 940 -865 960 -840
rect 940 -885 960 -865
rect 2095 -845 2140 -825
rect 1095 -1195 1115 -925
rect 1295 -1195 1315 -925
rect 1495 -1195 1515 -925
rect 1695 -1195 1715 -925
rect 1895 -1195 1915 -925
rect 2095 -1195 2115 -925
rect 1195 -1315 1240 -1295
rect 70 -1375 115 -1355
rect 70 -1490 90 -1445
rect 195 -1440 215 -1395
rect 295 -1440 315 -1395
rect 495 -1440 515 -1395
rect 695 -1440 715 -1395
rect 895 -1440 915 -1395
rect 1095 -1440 1115 -1395
rect 1145 -1440 1165 -1395
rect 1195 -1440 1215 -1395
rect 1395 -1440 1415 -1395
rect 1595 -1440 1615 -1395
rect 1795 -1440 1815 -1395
rect 1995 -1440 2015 -1395
rect 2095 -1440 2115 -1395
<< metal1 >>
rect 180 -200 2130 -190
rect 180 -245 195 -200
rect 215 -245 295 -200
rect 315 -245 495 -200
rect 515 -245 695 -200
rect 715 -245 895 -200
rect 915 -245 1095 -200
rect 1115 -245 1145 -200
rect 1165 -245 1195 -200
rect 1215 -245 1395 -200
rect 1415 -245 1595 -200
rect 1615 -245 1795 -200
rect 1815 -245 1995 -200
rect 2015 -245 2095 -200
rect 2115 -245 2130 -200
rect 180 -255 2130 -245
rect 285 -425 325 -255
rect 2085 -425 2125 -255
rect 60 -435 2125 -425
rect 60 -705 95 -435
rect 115 -705 295 -435
rect 315 -705 495 -435
rect 515 -705 695 -435
rect 715 -705 895 -435
rect 915 -705 1095 -435
rect 1115 -705 2095 -435
rect 2115 -705 2125 -435
rect 60 -715 2125 -705
rect 2085 -825 2150 -815
rect 2085 -830 2095 -825
rect 930 -840 2095 -830
rect 930 -885 940 -840
rect 960 -845 2095 -840
rect 2140 -845 2150 -825
rect 960 -855 2150 -845
rect 960 -885 970 -855
rect 930 -895 970 -885
rect 60 -925 2125 -915
rect 60 -1195 95 -925
rect 115 -1195 1095 -925
rect 1115 -1195 1295 -925
rect 1315 -1195 1495 -925
rect 1515 -1195 1695 -925
rect 1715 -1195 1895 -925
rect 1915 -1195 2095 -925
rect 2115 -1195 2125 -925
rect 60 -1205 2125 -1195
rect 140 -1295 1250 -1285
rect 140 -1315 1195 -1295
rect 1240 -1315 1250 -1295
rect 140 -1325 1250 -1315
rect 60 -1355 125 -1345
rect 60 -1375 70 -1355
rect 115 -1375 125 -1355
rect 60 -1385 125 -1375
rect 140 -1435 165 -1325
rect 1385 -1385 1425 -1205
rect 2085 -1385 2125 -1205
rect 60 -1445 165 -1435
rect 60 -1490 70 -1445
rect 90 -1490 165 -1445
rect 180 -1395 2130 -1385
rect 180 -1440 195 -1395
rect 215 -1440 295 -1395
rect 315 -1440 495 -1395
rect 515 -1440 695 -1395
rect 715 -1440 895 -1395
rect 915 -1440 1095 -1395
rect 1115 -1440 1145 -1395
rect 1165 -1440 1195 -1395
rect 1215 -1440 1395 -1395
rect 1415 -1440 1595 -1395
rect 1615 -1440 1795 -1395
rect 1815 -1440 1995 -1395
rect 2015 -1440 2095 -1395
rect 2115 -1440 2130 -1395
rect 180 -1450 2130 -1440
rect 60 -1500 165 -1490
<< labels >>
rlabel metal1 60 -1055 60 -1055 7 VP
port 1 w
rlabel metal1 60 -570 60 -570 7 VN
port 2 w
rlabel locali 60 -340 60 -340 7 I1p
port 3 w
rlabel locali 60 -745 60 -745 7 Vbn
port 4 w
rlabel locali 60 -1365 60 -1365 7 I1n
port 5 w
rlabel locali 60 -1465 60 -1465 7 Vbp
port 6 w
rlabel locali 2150 -745 2150 -745 3 Vcn
port 8 e
rlabel locali 2150 -835 2150 -835 3 Vcp
port 7 e
<< end >>
